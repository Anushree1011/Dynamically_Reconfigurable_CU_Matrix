library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.custom_pack.all;
use std.env.finish;
entity final_tb is
end final_tb;
architecture Behavioral of final_tb is
constant d_w_c: integer := 4;
signal input1,input2: arr_1d(0 to 3)(d_w_c-1 downto 0);
signal Sel: arr_2d(0 to 3)(0 to 3)(4 downto 0);
signal mux_sel: arr_2d(0 to 3)(0 to 7)(1 downto 0);
signal cu_Output: arr_2d(0 to 3)(0 to 3)(d_w_c-1 downto 0);
signal clk: std_logic:= '0';
signal w_en_ina, w_en_inb, w_en_in, w_en_out :arr_2d_b(0 to 3)(0 to 3);
signal final_output: arr_1d(0 to 3)(d_w_c - 1 downto 0);
begin
dut: entity work.final(Behavioral)
generic map(d_w => d_w_c)
port map(
input1 => input1, input2 => input2, mux_sel => mux_sel, Sel => Sel, cu_Output => cu_Output, final_output => final_output, clk => clk, w_en_in => w_en_in, w_en_out => w_en_out, w_en_ina => w_en_ina, w_en_inb => w_en_inb);
clk <= not clk after 5 ns;
process
begin

--RUN 1
input1(0)<="1010";input2(0)<="0100";input1(1)<="1101";input2(1)<="1011";input1(2)<="1010";input2(2)<="1010";input1(3)<="1100";input2(3)<="1010";
mux_sel(0)(0)<="00";mux_sel(0)(1)<="00";mux_sel(0)(2)<="01";mux_sel(0)(3)<="00";mux_sel(0)(4)<="01";mux_sel(0)(5)<="01";mux_sel(0)(6)<="00";mux_sel(0)(7)<="01";
Sel(0)(0)<="00111";Sel(0)(1)<="01000";Sel(0)(2)<="00110";Sel(0)(3)<="10011";
w_en_ina(0)(0) <= '1';
w_en_inb(0)(0) <= '1'; 
w_en_in(0)(0) <= '1'; wait for 10ns;
w_en_ina(0)(0) <= '0'; 
w_en_inb(0)(0) <= '0'; 
w_en_in(0)(0) <= '0'; 
w_en_out(0)(0) <= '1'; wait for 20 ns;
w_en_out(0)(0) <= '0'; wait for 10 ns;
w_en_ina(0)(1) <= '1'; 
w_en_inb(0)(1) <= '1';
w_en_in(0)(1) <= '1'; wait for 10ns;
w_en_ina(0)(1) <= '0';
w_en_inb(0)(1) <= '0';
w_en_in(0)(1) <= '0';
w_en_out(0)(1) <= '1';wait for 20 ns;
w_en_out(0)(1) <= '0'; wait for 10 ns;
w_en_ina(0)(2) <= '1'; 
w_en_inb(0)(2) <= '1'; 
w_en_in(0)(2) <= '1'; wait for 20 ns;
w_en_ina(0)(2) <= '0'; 
w_en_inb(0)(2) <= '0'; 
w_en_in(0)(2) <= '0'; 
w_en_out(0)(2) <= '1'; wait for 20 ns;
w_en_out(0)(2) <= '0'; wait for 10 ns;
w_en_ina(0)(3) <= '1';
w_en_inb(0)(3) <= '1';
w_en_in(0)(3) <= '1';wait for 10 ns;
w_en_ina(0)(3) <= '0'; 
w_en_inb(0)(3) <= '0'; 
w_en_in(0)(3) <= '0'; 
w_en_out(0)(3) <= '1';wait for 20 ns;
w_en_out(0)(3) <= '0'; wait for 10 ns;
mux_sel(1)(0)<="00";mux_sel(1)(1)<="00";mux_sel(1)(2)<="01";mux_sel(1)(3)<="00";mux_sel(1)(4)<="01";mux_sel(1)(5)<="00";mux_sel(1)(6)<="01";mux_sel(1)(7)<="01";
Sel(1)(0)<="10010";Sel(1)(1)<="10100";Sel(1)(2)<="01110";Sel(1)(3)<="01100";
w_en_ina(1)(0) <= '1';
w_en_inb(1)(0) <= '1';
w_en_in(1)(0) <= '1'; wait for 10ns;
w_en_ina(1)(0) <= '0';
w_en_inb(1)(0) <= '0'; 
w_en_in(1)(0) <= '0'; 
w_en_out(1)(0) <= '1';wait for 20 ns;
w_en_out(1)(0) <= '0';wait for 10 ns;
w_en_ina(1)(1) <= '1';
w_en_inb(1)(1) <= '1'; 
w_en_in(1)(1) <= '1'; wait for 10ns;
w_en_ina(1)(1) <= '0';
w_en_inb(1)(1) <= '0';
w_en_in(1)(1) <= '0';
w_en_out(1)(1) <= '1'; wait for 20ns;
w_en_out(1)(1) <= '0'; wait for 10ns;
w_en_ina(1)(2) <= '1'; 
w_en_inb(1)(2) <= '1'; 
w_en_in(1)(2) <= '1'; wait for 10ns;
w_en_ina(1)(2) <= '0'; 
w_en_inb(1)(2) <= '0'; 
w_en_in(1)(2) <= '0'; 
w_en_out(1)(2) <= '1';wait for 20ns;
w_en_out(1)(2) <= '0'; wait for 10ns;
w_en_ina(1)(3) <= '1';
w_en_inb(1)(3) <= '1';
w_en_in(1)(3) <= '1';wait for 10 ns;
w_en_ina(1)(3) <= '0'; 
w_en_inb(1)(3) <= '0';
w_en_in(1)(3) <= '0'; 
w_en_out(1)(3) <= '1';wait for 20 ns;
w_en_out(1)(3) <= '0'; wait for 10 ns;
mux_sel(2)(0)<="00";mux_sel(2)(1)<="01";mux_sel(2)(2)<="10";mux_sel(2)(3)<="00";mux_sel(2)(4)<="10";mux_sel(2)(5)<="01";mux_sel(2)(6)<="01";mux_sel(2)(7)<="00";
Sel(2)(0)<="00101";Sel(2)(1)<="10101";Sel(2)(2)<="00011";Sel(2)(3)<="00001";
w_en_ina(2)(0) <= '1'; 
w_en_inb(2)(0) <= '1';
w_en_in(2)(0) <= '1'; wait for 10ns;
w_en_ina(2)(0) <= '0'; 
w_en_inb(2)(0) <= '0'; 
w_en_in(2)(0) <= '0'; 
w_en_out(2)(0) <= '1';wait for 20ns;
w_en_out(2)(0) <= '0';wait for 10ns;
w_en_ina(2)(1) <= '1'; 
w_en_inb(2)(1) <= '1'; 
w_en_in(2)(1) <= '1'; wait for 10ns;
w_en_ina(2)(1) <= '0'; 
w_en_inb(2)(1) <= '0'; 
w_en_in(2)(1) <= '0'; 
w_en_out(2)(1) <= '1';wait for 20ns;
w_en_out(2)(1) <= '0';wait for 10ns;
w_en_ina(2)(2) <= '1'; 
w_en_inb(2)(2) <= '1'; 
w_en_in(2)(2) <= '1'; wait for 10ns;
w_en_ina(2)(2) <= '0'; 
w_en_inb(2)(2) <= '0'; 
w_en_in(2)(2) <= '0'; 
w_en_out(2)(2) <= '1'; wait for 20ns;
w_en_out(2)(2) <= '0'; wait for 10ns;
w_en_ina(2)(3) <= '1';
w_en_inb(2)(3) <= '1';
w_en_in(2)(3) <= '1';wait for 10 ns;
w_en_ina(2)(3) <= '0'; 
w_en_inb(2)(3) <= '0'; 
w_en_in(2)(3) <= '0'; 
w_en_out(2)(3) <= '1';wait for 20 ns;
w_en_out(2)(3) <= '0'; wait for 10 ns;
mux_sel(3)(0)<="01";mux_sel(3)(1)<="00";mux_sel(3)(2)<="01";mux_sel(3)(3)<="10";mux_sel(3)(4)<="00";mux_sel(3)(5)<="01";mux_sel(3)(6)<="10";mux_sel(3)(7)<="00";
Sel(3)(0)<="10011";Sel(3)(1)<="01101";Sel(3)(2)<="01000";Sel(3)(3)<="00010";
w_en_ina(3)(0) <= '1';
w_en_inb(3)(0) <= '1';
w_en_in(3)(0) <= '1';wait for 10ns;
w_en_ina(3)(0) <= '0';
w_en_inb(3)(0) <= '0';
w_en_in(3)(0) <= '0'; 
w_en_out(3)(0) <= '1';wait for 20ns;
w_en_out(3)(0) <= '0';wait for 10ns;
w_en_ina(3)(1) <= '1'; 
w_en_inb(3)(1) <= '1'; 
w_en_in(3)(1) <= '1'; wait for 10 ns;
w_en_ina(3)(1) <= '0'; 
w_en_inb(3)(1) <= '0'; 
w_en_in(3)(1) <= '0'; 
w_en_out(3)(1) <= '1'; wait for 20 ns; 
w_en_out(3)(1) <= '0'; wait for 10 ns;
w_en_ina(3)(2) <= '1'; 
w_en_inb(3)(2) <= '1'; 
w_en_in(3)(2) <= '1'; wait for 10 ns;
w_en_ina(3)(2) <= '0'; 
w_en_inb(3)(2) <= '0'; 
w_en_in(3)(2) <= '0'; 
w_en_out(3)(2) <= '1'; wait for 20 ns;
w_en_out(3)(2) <= '0'; wait for 10 ns;
w_en_ina(3)(3) <= '1';
w_en_inb(3)(3) <= '1';
w_en_in(3)(3) <= '1';wait for 10 ns;
w_en_ina(3)(3) <= '0'; 
w_en_inb(3)(3) <= '0'; 
w_en_in(3)(3) <= '0'; 
w_en_out(3)(3) <= '1';wait for 20 ns;
w_en_out(3)(3) <= '0'; wait for 10 ns;

--Run 2

mux_sel(0)(0)<="01";mux_sel(0)(1)<="01";mux_sel(0)(2)<="01";mux_sel(0)(3)<="10";mux_sel(0)(4)<="10";mux_sel(0)(5)<="01";mux_sel(0)(6)<="10";mux_sel(0)(7)<="01";
Sel(0)(0)<="00100";Sel(0)(1)<="00101";Sel(0)(2)<="00011";Sel(0)(3)<="01000";
w_en_ina(0)(0) <= '1';
w_en_inb(0)(0) <= '1'; 
w_en_in(0)(0) <= '1'; wait for 10ns;
w_en_ina(0)(0) <= '0'; 
w_en_inb(0)(0) <= '0'; 
w_en_in(0)(0) <= '0'; 
w_en_out(0)(0) <= '1'; wait for 20 ns;
w_en_out(0)(0) <= '0'; wait for 10 ns;
w_en_ina(0)(1) <= '1'; 
w_en_inb(0)(1) <= '1';
w_en_in(0)(1) <= '1'; wait for 10ns;
w_en_ina(0)(1) <= '0';
w_en_inb(0)(1) <= '0';
w_en_in(0)(1) <= '0';
w_en_out(0)(1) <= '1';wait for 20 ns;
w_en_out(0)(1) <= '0'; wait for 10 ns;
w_en_ina(0)(2) <= '1'; 
w_en_inb(0)(2) <= '1'; 
w_en_in(0)(2) <= '1'; wait for 20 ns;
w_en_ina(0)(2) <= '0'; 
w_en_inb(0)(2) <= '0'; 
w_en_in(0)(2) <= '0'; 
w_en_out(0)(2) <= '1'; wait for 20 ns;
w_en_out(0)(2) <= '0'; wait for 10 ns;
w_en_ina(0)(3) <= '1';
w_en_inb(0)(3) <= '1';
w_en_in(0)(3) <= '1';wait for 10 ns;
w_en_ina(0)(3) <= '0'; 
w_en_inb(0)(3) <= '0'; 
w_en_in(0)(3) <= '0'; 
w_en_out(0)(3) <= '1';wait for 20 ns;
w_en_out(0)(3) <= '0'; wait for 10 ns;
mux_sel(1)(0)<="00";mux_sel(1)(1)<="00";mux_sel(1)(2)<="01";mux_sel(1)(3)<="00";mux_sel(1)(4)<="01";mux_sel(1)(5)<="00";mux_sel(1)(6)<="01";mux_sel(1)(7)<="00";
Sel(1)(0)<="00111";Sel(1)(1)<="01100";Sel(1)(2)<="00110";Sel(1)(3)<="01110";
w_en_ina(1)(0) <= '1';
w_en_inb(1)(0) <= '1';
w_en_in(1)(0) <= '1'; wait for 10ns;
w_en_ina(1)(0) <= '0';
w_en_inb(1)(0) <= '0'; 
w_en_in(1)(0) <= '0'; 
w_en_out(1)(0) <= '1';wait for 20 ns;
w_en_out(1)(0) <= '0';wait for 10 ns;
w_en_ina(1)(1) <= '1';
w_en_inb(1)(1) <= '1'; 
w_en_in(1)(1) <= '1'; wait for 10ns;
w_en_ina(1)(1) <= '0';
w_en_inb(1)(1) <= '0';
w_en_in(1)(1) <= '0';
w_en_out(1)(1) <= '1'; wait for 20ns;
w_en_out(1)(1) <= '0'; wait for 10ns;
w_en_ina(1)(2) <= '1'; 
w_en_inb(1)(2) <= '1'; 
w_en_in(1)(2) <= '1'; wait for 10ns;
w_en_ina(1)(2) <= '0'; 
w_en_inb(1)(2) <= '0'; 
w_en_in(1)(2) <= '0'; 
w_en_out(1)(2) <= '1';wait for 20ns;
w_en_out(1)(2) <= '0'; wait for 10ns;
w_en_ina(1)(3) <= '1';
w_en_inb(1)(3) <= '1';
w_en_in(1)(3) <= '1';wait for 10 ns;
w_en_ina(1)(3) <= '0'; 
w_en_inb(1)(3) <= '0';
w_en_in(1)(3) <= '0'; 
w_en_out(1)(3) <= '1';wait for 20 ns;
w_en_out(1)(3) <= '0'; wait for 10 ns;
mux_sel(2)(0)<="01";mux_sel(2)(1)<="00";mux_sel(2)(2)<="10";mux_sel(2)(3)<="00";mux_sel(2)(4)<="00";mux_sel(2)(5)<="01";mux_sel(2)(6)<="01";mux_sel(2)(7)<="00";
Sel(2)(0)<="10010";Sel(2)(1)<="01011";Sel(2)(2)<="01000";Sel(2)(3)<="00001";
w_en_ina(2)(0) <= '1'; 
w_en_inb(2)(0) <= '1';
w_en_in(2)(0) <= '1'; wait for 10ns;
w_en_ina(2)(0) <= '0'; 
w_en_inb(2)(0) <= '0'; 
w_en_in(2)(0) <= '0'; 
w_en_out(2)(0) <= '1';wait for 20ns;
w_en_out(2)(0) <= '0';wait for 10ns;
w_en_ina(2)(1) <= '1'; 
w_en_inb(2)(1) <= '1'; 
w_en_in(2)(1) <= '1'; wait for 10ns;
w_en_ina(2)(1) <= '0'; 
w_en_inb(2)(1) <= '0'; 
w_en_in(2)(1) <= '0'; 
w_en_out(2)(1) <= '1';wait for 20ns;
w_en_out(2)(1) <= '0';wait for 10ns;
w_en_ina(2)(2) <= '1'; 
w_en_inb(2)(2) <= '1'; 
w_en_in(2)(2) <= '1'; wait for 10ns;
w_en_ina(2)(2) <= '0'; 
w_en_inb(2)(2) <= '0'; 
w_en_in(2)(2) <= '0'; 
w_en_out(2)(2) <= '1'; wait for 20ns;
w_en_out(2)(2) <= '0'; wait for 10ns;
w_en_ina(2)(3) <= '1';
w_en_inb(2)(3) <= '1';
w_en_in(2)(3) <= '1';wait for 10 ns;
w_en_ina(2)(3) <= '0'; 
w_en_inb(2)(3) <= '0'; 
w_en_in(2)(3) <= '0'; 
w_en_out(2)(3) <= '1';wait for 20 ns;
w_en_out(2)(3) <= '0'; wait for 10 ns;
mux_sel(3)(0)<="00";mux_sel(3)(1)<="01";mux_sel(3)(2)<="00";mux_sel(3)(3)<="10";mux_sel(3)(4)<="00";mux_sel(3)(5)<="10";mux_sel(3)(6)<="01";mux_sel(3)(7)<="10";
Sel(3)(0)<="01001";Sel(3)(1)<="10101";Sel(3)(2)<="10001";Sel(3)(3)<="10100";
w_en_ina(3)(0) <= '1';
w_en_inb(3)(0) <= '1';
w_en_in(3)(0) <= '1';wait for 10ns;
w_en_ina(3)(0) <= '0';
w_en_inb(3)(0) <= '0';
w_en_in(3)(0) <= '0'; 
w_en_out(3)(0) <= '1';wait for 20ns;
w_en_out(3)(0) <= '0';wait for 10ns;
w_en_ina(3)(1) <= '1'; 
w_en_inb(3)(1) <= '1'; 
w_en_in(3)(1) <= '1'; wait for 10 ns;
w_en_ina(3)(1) <= '0'; 
w_en_inb(3)(1) <= '0'; 
w_en_in(3)(1) <= '0'; 
w_en_out(3)(1) <= '1'; wait for 20 ns; 
w_en_out(3)(1) <= '0'; wait for 10 ns;
w_en_ina(3)(2) <= '1'; 
w_en_inb(3)(2) <= '1'; 
w_en_in(3)(2) <= '1'; wait for 10 ns;
w_en_ina(3)(2) <= '0'; 
w_en_inb(3)(2) <= '0'; 
w_en_in(3)(2) <= '0'; 
w_en_out(3)(2) <= '1'; wait for 20 ns;
w_en_out(3)(2) <= '0'; wait for 10 ns;
w_en_ina(3)(3) <= '1';
w_en_inb(3)(3) <= '1';
w_en_in(3)(3) <= '1';wait for 10 ns;
w_en_ina(3)(3) <= '0'; 
w_en_inb(3)(3) <= '0'; 
w_en_in(3)(3) <= '0'; 
w_en_out(3)(3) <= '1';wait for 20 ns;
w_en_out(3)(3) <= '0'; wait for 20 ns;

finish;
end process;
end Behavioral;

